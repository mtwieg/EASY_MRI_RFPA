** Profile: "SCHEMATIC1-TransientAnalysis"  [ C:\Users\a0232073\Downloads\LM7171\lm7171-pspicefiles\schematic1\transientanalysis.sim ] 

** Creating circuit file "TransientAnalysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../LM7171.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 0.1e-9 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 N([VOUT])
.INC "..\SCHEMATIC1.net" 


.END
