*Feb 19, 2010 *Doc. ID: 90199, Rev. A *File Name: part irf630_sihf630_PS.txt and part irf630_sihf630_PS.spi *This document is intended as a SPICE modeling guideline and does not *constitute a commercial product datasheet. Designers should refer to the *appropriate data sheet of the same number for guaranteed specification *limits. .SUBCKT irf630 1 2 3 ************************************** * Model Generated by MODPEX * *Copyright(c) Symmetry Design Systems* * All Rights Reserved * * UNPUBLISHED LICENSED SOFTWARE * * Contains Proprietary Information * * Which is The Property of * * SYMMETRY OR ITS LICENSORS * *Commercial Use or Resale Restricted * * by Symmetry License Agreement * ************************************** * Model generated on Jun 25, 96 * Model format: SPICE3 * Symmetry POWER MOS Model (Version 1.0) * External Node Designations * Node 1 -> Drain * Node 2 -> Gate * Node 3 -> Source M1 9 7 8 8 MM L=100u W=100u * Default values used in MM: * The voltage-dependent capacitances are * not included. Other default values are: * RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0 .MODEL MM NMOS LEVEL=1 IS=1e-32 +VTO=3.90614 LAMBDA=0 KP=2.70091 +CGSO=7.25845e-06 CGDO=1e-11 RS 8 3 0.0001 D1 3 1 MD .MODEL MD D IS=2.59955e-15 RS=0.0232241 N=0.818263 BV=200 +IBV=0.00025 EG=1 XTI=2.54918 TT=0 +CJO=6.35847e-10 VJ=5 M=0.772431 FC=0.5 RDS 3 1 8e+06 RD 9 1 0.169992 RG 2 7 4.09017 D2 4 5 MD1 * Default values used in MD1: * RS=0 EG=1.11 XTI=3.0 TT=0 * BV=infinite IBV=1mA .MODEL MD1 D IS=1e-32 N=50 +CJO=1.28188e-09 VJ=1.20026 M=0.9 FC=1e-08 D3 0 5 MD2 * Default values used in MD2: * EG=1.11 XTI=3.0 TT=0 CJO=0 * BV=infinite IBV=1mA .MODEL MD2 D IS=1e-10 N=0.413904 RS=3e-06 RL 5 10 1 FI2 7 9 VFI2 -1 VFI2 4 0 0 EV16 10 0 9 7 1 CAP 11 10 1.2819e-09 FI1 7 9 VFI1 -1 VFI1 11 6 0 RCAP 6 10 1 D4 0 6 MD3 * Default values used in MD3: * EG=1.11 XTI=3.0 TT=0 CJO=0 * RS=0 BV=infinite IBV=1mA .MODEL MD3 D IS=1e-10 N=0.413904 .ENDS